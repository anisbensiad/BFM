package dual_protocol_pkg;
    // Memory load structure
    typedef struct {
        string memory_path;
        string data_file_path;
    } mem_load_t;
endpackage
